module core();
endmodule
